//p19
library ieee;
use ieee.std_logic_1164.all;

entity and_gate is 
   port(a1,a2: in std_logic;
        b1:    out std_logic
       );
 end and_gate;

architecture behav of and_gate is
  begin 
     b1<= a1 and a2;
end behav;

//p20
library ieee;
use ieee.std_logic_1164.all;

entity or_gate is 
  port(a1,a2: in std_logic;
       b1:    out std_logic
      );
end or_gate;

architecture behav of or_gate is 
   begin 
     b1<=a1 or a2;
end behav;

//p26
library ieee;
use ieee.std_logic_1164.all;

entity COUNTER is 
  port(clk: in std_logic;
       rs:  in std_logic;
       count_out: out std_logic_vector(2 downto 0)
      );
end COUNTER;

architecture behav of COUNTER is 
   signal next_counter: std_logic_vector(2 downto 0);
   begin 
      process(rs,clk)
         begin 
            if rs='0' then next_counter <="000";
              elsif (clk'event and clk='1') then
                  case next_counter is 
                     when "000" => next_counter<="001";
                     when "001" => next_counter<="011";
                     when "011" => next_counter<="111";
                     when "111" => next_counter<="110";
                     when "110" => next_counter<="100";
                     when "100" => next_counter<="000";
                     when others => next_counter<="XXX";
                  end case;
            end if;
            count_out <= next_counter;
      end process;
 end behav;

//p34
-- megafunction wizard: %LPM_RAM_DP%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: memory.vhd
-- Megafunction Name(s):
-- 			altsyncram
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 5.1 Build 176 10/26/2005 SJ Full Version
-- ************************************************************
LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY memory IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		rdaddress		: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		wraddress		: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		wren		: IN STD_LOGIC  := '1';
		q		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END memory;


ARCHITECTURE SYN OF memory IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);



	COMPONENT altsyncram
	GENERIC (
		address_reg_b		: STRING;
		clock_enable_input_a		: STRING;
		clock_enable_input_b		: STRING;
		clock_enable_output_b		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		numwords_a		: NATURAL;
		numwords_b		: NATURAL;
		operation_mode		: STRING;
		outdata_aclr_b		: STRING;
		outdata_reg_b		: STRING;
		power_up_uninitialized		: STRING;
		read_during_write_mode_mixed_ports		: STRING;
		widthad_a		: NATURAL;
		widthad_b		: NATURAL;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_byteena_a		: NATURAL
	);
	PORT (
			wren_a	: IN STD_LOGIC ;
			clock0	: IN STD_LOGIC ;
			address_a	: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
			address_b	: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
			q_b	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			data_a	: IN STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	q    <= sub_wire0(15 DOWNTO 0);

	altsyncram_component : altsyncram
	GENERIC MAP (
		address_reg_b => "CLOCK0",
		clock_enable_input_a => "BYPASS",
		clock_enable_input_b => "BYPASS",
		clock_enable_output_b => "BYPASS",
		intended_device_family => "Cyclone II",
		lpm_type => "altsyncram",
		numwords_a => 64,
		numwords_b => 64,
		operation_mode => "DUAL_PORT",
		outdata_aclr_b => "NONE",
		outdata_reg_b => "UNREGISTERED",
		power_up_uninitialized => "FALSE",
		read_during_write_mode_mixed_ports => "DONT_CARE",
		widthad_a => 6,
		widthad_b => 6,
		width_a => 16,
		width_b => 16,
		width_byteena_a => 1
	)
	PORT MAP (
		wren_a => wren,
		clock0 => clock,
		address_a => wraddress,
		address_b => rdaddress,
		data_a => data,
		q_b => sub_wire0
	);
END SYN;
    
//p51
library ieee;
use ieee.std_logic_1164.all;

entity register_16 is port
   (reset:   in std_logic;
    d_input: in std_logic_vector(15 downto 0);
    clk:     in std_logic;
    write:   in std_logic;
    sel:     in std_logic;
    q_output: out std_logic_vector(15 downto 0)
   );
end register_16;

architecture a of register_16 is 
   begin 
      process(reset,clk)
         begin      
           if reset='0' then 
              q_output<=x"0000";
            elsif(clk'event and clk='1') then
               if sel='1' and write='1' then 
                  q_output<=d_input;
         end if;
      end if;
   end process;
end a;
  
 （2）设计实体decoder2_to_4
library ieee;
use ieee.std_logic_1164.all;

entity decoder2_to_4 is 
  port(sel: in std_logic_vector(1 downto 0);
       sel00: out std_logic;
       sel01: out std_logic;
       sel02: out std_logic;
       sel03: out std_logic
      );
end decoder2_to_4;

architecture behavioral of decoder2_to_4 is 
   begin 
     sel00<=(not sel(1)) and (not sel(0));
     sel01<=(not sel(1)) and sel(0);
     sel02<= sel(1) and (not sel(0));
     sel03<= sel(1) and sel(0);
   end behavioral;

（3）设计实体mux4_to_1
ibrary ieee;
use ieee.std_logic_1164.all;

entity mux4_to_1 is 
   port(input0,input1,input2,input3: in std_logic_vector(15 downto 0);
        sel:  in std_logic_vector(1 downto 0);
        out_put: out std_logic_vector(15 downto 0));
end mux4_to_1;

architecture behavioral of mux4_to_1 is 
  begin 
    mux: process(sel, input0,input1,input2,input3)
         begin 
            case sel is
                when "00" => out_put<= input0;
                when "01" => out_put<= input1;
                when "10" => out_put<= input2;
                when "11" => out_put<= input3;
            end case;
    end process;
end behavioral;

（4）高层设计实体regfile
library ieee;
use ieee.std_logic_1164.all;

entity regfile is
  port(DR: in std_logic_vector(1 downto 0);
       SR: in std_logic_vector(1 downto 0);
       reset:   in std_logic;
       DRWr:    in std_logic;
       clk:     in std_logic;
       d_input: in std_logic_vector(15 downto 0);
       DR_data: out std_logic_vector(15 downto 0);
       SR_data: out std_logic_vector(15 downto 0)
      );
end regfile;

architecture struct of regfile is 
   component register_16
      port(reset,clk,write,sel: in std_logic;
           d_input: in std_logic_vector(15 downto 0);
           q_output: out std_logic_vector(15 downto 0)
           );
   end component;

   component decoder2_to_4
      port(sel: in std_logic_vector(1 downto 0);
           sel00,sel01,sel02,sel03: out std_logic
           );
   end component;

    component mux4_to_1
      port(input0,input1,input2,input3: in std_logic_vector(15 downto 0);
           sel:     in std_logic_vector(1 downto 0);
           out_put: out std_logic_vector(15 downto 0)
           );
   end component;

       signal reg00,reg01,reg02,reg03: std_logic_vector(15 downto 0);
       signal sel00,sel01,sel02,sel03: std_logic;

   begin
     Areg00:register_16 port map(
             reset   => reset,
             d_input => d_input,
             clk     => clk,
             write   => DRWr,
             sel     => sel00,
             q_output=> reg00
            );
     Areg01:register_16 port map(
             reset   => reset,
             d_input => d_input,
             clk     => clk,
             write   => DRWr,
             sel     => sel01,
             q_output=> reg01
            );
      Areg02:register_16 port map(
             reset   => reset,
             d_input => d_input,
             clk     => clk,
             write   => DRWr,
             sel     => sel02,
             q_output=> reg02
            );
      Areg03:register_16 port map(
             reset   => reset,
             d_input => d_input,
             clk     => clk,
             write   => DRWr,
             sel     => sel03,
             q_output=> reg03
            );
       decoder: decoder2_to_4 port map(
             sel     => DR,
             sel00   => sel00,
             sel01   => sel01,
             sel02   => sel02,
             sel03   => sel03
           );
       mux1:  mux4_to_1 port map(
             input0 => reg00,
             input1 => reg01,
             input2 => reg02,
             input3 => reg03,
             sel    => DR,
             out_put =>DR_data
           );
        mux2:  mux4_to_1 port map(
             input0 => reg00,
             input1 => reg01,
             input2 => reg02,
             input3 => reg03,
             sel    => SR,
             out_put =>SR_data
           );
end struct;

//p60
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity alu is
port(cin:in std_logic;
     alu_a,alu_b:in std_logic_vector(15 downto 0);
     alu_func:in std_logic_vector(2 downto 0);
     alu_out:out std_logic_vector(15 downto 0);
     c,z,v,s:out std_logic);
end alu;

architecture behave of alu is
begin
	process(alu_a,alu_b,cin,alu_func)
	variable temp1,temp2,temp3 : std_logic_vector(15 downto 0) ;
	begin
		temp1 := "000000000000000"&cin;
		case alu_func is
			when "000"=>
			temp2 := alu_b+alu_a+temp1;
			when "001"=>
			temp2 := alu_b-alu_a-temp1;
			when "010"=>
			temp2 := alu_a and alu_b;
			when "011"=>
			temp2 := alu_a or alu_b;
			when "100"=>
			temp2 := alu_a xor alu_b;
			when "101"=>
			temp2(0) := '0';
			for I in 15 downto 1 loop
			temp2(I) := alu_b(I-1);
			end loop;
			when "110"=>
			temp2(15) := '0';
			for I in 14 downto 0 loop
			temp2(I) := alu_b(I+1);
			end loop;
			when others=>
			temp2 := "0000000000000000";
		end case;
		alu_out <= temp2;
		if temp2 = "0000000000000000" then z<='1';
		else z<='0';
		end if;
		if temp2(15) = '1' then s<='1';
		else s<='0';
		end if;
		case alu_func is
			when "000" | "001"=>
			if (alu_a(15)= '1' and alu_b(15)= '1' and temp2(15) = '0') or
			   (alu_a(15)= '0' and alu_b(15)= '0' and temp2(15) = '1') then
			v<='1';
			else v<='0';
			end if;
			when others=>
			v<='0';
		end case;
		case alu_func is
			when "000"=>
			temp3 := "1111111111111111"-alu_b-temp1;
			if temp3<alu_a then
			c<='1';
			else c<='0';
			end if;
			when "001"=>
			if alu_b<alu_a then
			c<='1';
			else c<='0';
			end if;
			when "101"=>
			c <= alu_b(15);
			when "110"=>
			c <= alu_b(0);
			when others=>
			c<='0';
		end case;
	end process;
end behave;

//p62
library ieee;
use ieee.std_logic_1164.all;

entity reg is
	port(d:            in std_logic_vector(15 downto 0);
	     clk,reset,en: in std_logic;
	     q:out std_logic_vector(15 downto 0));
end reg;

architecture behave of reg is
begin
	process(clk,reset,en)
	begin
		if reset = '0' then            
          q <= "0000000000000000";
        elsif clk'event and clk = '1' then
          if en = '1' then
			q <= d;
		  end if;
        end if;
	end process;
end behave;

//p70
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity alu is
port(cin:in std_logic;
     alu_a,alu_b:in std_logic_vector(15 downto 0);
     alu_func:in std_logic_vector(2 downto 0);
     alu_out:out std_logic_vector(15 downto 0);
     c,z,v,s:out std_logic);
end alu;

architecture behave of alu is
begin
	process(alu_a,alu_b,cin,alu_func)
	variable temp1,temp2,temp3 : std_logic_vector(15 downto 0) ;
	begin
		temp1 := "000000000000000"&cin;
		case alu_func is
			when "000"=>
			temp2 := alu_b+alu_a+temp1;
			when "001"=>
			temp2 := alu_b-alu_a-temp1;
			when "010"=>
			temp2 := alu_a and alu_b;
			when "011"=>
			temp2 := alu_a or alu_b;
			when "100"=>
			temp2 := alu_a xor alu_b;
			when "101"=>
			temp2(0) := '0';
			for I in 15 downto 1 loop
			temp2(I) := alu_b(I-1);
			end loop;
			when "110"=>
			temp2(15) := '0';
			for I in 14 downto 0 loop
			temp2(I) := alu_b(I+1);
			end loop;
			when others=>
			temp2 := "0000000000000000";
		end case;
		alu_out <= temp2;
		if temp2 = "0000000000000000" then z<='1';
		else z<='0';
		end if;
		if temp2(15) = '1' then s<='1';
		else s<='0';
		end if;
		case alu_func is
			when "000" | "001"=>
			if (alu_a(15)= '1' and alu_b(15)= '1' and temp2(15) = '0') or
			   (alu_a(15)= '0' and alu_b(15)= '0' and temp2(15) = '1') then
			v<='1';
			else v<='0';
			end if;
			when others=>
			v<='0';
		end case;
		case alu_func is
			when "000"=>
			temp3 := "1111111111111111"-alu_b-temp1;
			if temp3<alu_a then
			c<='1';
			else c<='0';
			end if;
			when "001"=>
			if alu_b<alu_a then
			c<='1';
			else c<='0';
			end if;
			when "101"=>
			c <= alu_b(15);
			when "110"=>
			c <= alu_b(0);
			when others=>
			c<='0';
		end case;
	end process;
end behave;

//p71
library ieee;
use ieee.std_logic_1164.all;

entity reg is
	port
	(
		clr: 		in	std_logic;
		D:		 	in	std_logic_vector(15 downto 0);
		clock:		in	std_logic;
		write:		in	std_logic;
	    sel:		in	std_logic;
		Q:		 	out	std_logic_vector(15 downto 0)
	);
	
end reg;

architecture behav of reg is
begin
	process(clr,clock)
	begin
		if clr = '0' then
			Q <= x"0000"; 	
		elsif (clock'event and clock = '1') then
			if sel = '1' and write = '1' then
				Q <= D;
			end if;
		end if;
	end process;
end behav;

//p71
library ieee;
use ieee.std_logic_1164.all;

entity mux_4_to_1 is
port (
	input0,
	input1,
	input2,
	input3: 	in std_logic_vector(15 downto 0);
	sel: 		in std_logic_vector(1 downto 0);
	out_put: 	out std_logic_vector(15 downto 0));
end mux_4_to_1;

architecture behav of mux_4_to_1 is
begin
mux: process(sel, input0, input1, input2, input3)
begin
	case sel is 
		when "00" => 
			out_put <= input0;
		when "01" => 
			out_put <= input1;
		when "10" => 
			out_put <= input2;
		when "11" => 
			out_put <= input3;
	end case;
end process;
end behav;

//p74
Library ieee;
use ieee.std_logic_1164.all;

entity decoder_2_to_4 is	
    port (
		sel: 	in std_logic_vector(1 downto 0);
		sel00:  out std_logic;
		sel01:  out std_logic;
		sel02:  out std_logic;
		sel03:  out std_logic
		);
end decoder_2_to_4;

architecture behav of decoder_2_to_4 is
begin
	sel00	<=  (not sel(1)) and (not sel(0));
	sel01	<=  (not sel(1)) and sel(0) ;
	sel02	<=  sel(1) and (not sel(0)) ;
	sel03	<=  sel(1) and sel(0) ;
end behav;

//p74
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity regfile is
Port (  DR: 		in std_logic_vector(1 downto 0); 
		SR: 		in std_logic_vector(1 downto 0);   
		reset:  	in std_logic;
		DRWr:   	in std_logic;                           
		clk: 		in std_logic;	
		d_input: 	in  std_logic_vector(15 downto 0);
		DR_data:	out std_logic_vector(15 downto 0);        
		SR_data:  	out std_logic_vector(15 downto 0)   
	  );
end regfile;


architecture struct of regfile is
-- components
-- 16 bit Register for register file
component reg
port	(
		clr: 	in	std_logic;
		D: 		in	std_logic_vector(15 downto 0);
		clock: 	in	std_logic;
		write:  in	std_logic;
	    sel: 	in	std_logic;
		Q: 		out std_logic_vector(15 downto 0)
		);
end component;

-- 2 to 4 Decoder
component  decoder_2_to_4 
    port(
		sel: 	in  std_logic_vector(1 downto 0);
		sel00: 	out std_logic;
		sel01: 	out std_logic;
		sel02: 	out std_logic;
		sel03: 	out std_logic
		);
end component;

-- 4 to 1 line multiplexer
component mux_4_to_1
port (
	input0,
	input1,
	input2,
	input3:  in std_logic_vector(15 downto 0);
	sel:	 in std_logic_vector(1 downto 0);
	out_put: out std_logic_vector(15 downto 0));
end component;


signal reg00, reg01, reg02, reg03 
            :std_logic_vector(15 downto 0);
 
signal sel00 ,sel01 ,sel02 ,sel03
            : std_logic;

begin
Areg00: reg port map(
		clr			=>  reset,
		D			=>	d_input ,
		clock		=>	clk ,		
		write		=>	DRWr ,
	    sel			=>	sel00 ,	
		Q			=>  reg00
		);

Areg01: reg port map(
		clr			=>  reset,
		D			=>	d_input ,
		clock		=>	clk ,		
		write		=>	DRWr ,
	    sel			=>	sel01 ,	
		Q			=>  reg01	
		);

Areg02: reg port map(
		clr			=>  reset,
		D			=>  d_input ,
		clock		=>	clk ,		
		write		=>	DRWr ,
	    sel			=>	sel02 ,	
		Q			=>  reg02
		);

Areg03: reg port map(
		clr			=>  reset,
		D			=>	d_input ,
		clock		=>	clk ,		
		write		=>	DRWr ,
	    sel			=>	sel03 ,	
		Q			=>  reg03
		);

-- decoder
des_decoder: decoder_2_to_4 port map
		(
		sel 	=> DR,
    	sel00 	=> sel00 ,
		sel01 	=> sel01 ,
		sel02 	=> sel02 ,
		sel03 	=> sel03 
		);

mux1: mux_4_to_1 PORT MAP(
	Input0 => reg00 ,
    Input1 => reg01 ,
	Input2 => reg02 ,
	Input3 => reg03 ,
	sel => DR ,
	out_put => DR_data
	);
	
mux2: mux_4_to_1 PORT MAP(
	input0 	=> reg00 ,
    input1 	=> reg01 ,
	input2 	=> reg02 ,
	input3 	=> reg03 ,
	sel 	=> SR ,
	out_put => SR_data
	);

end struct;














